//commit 4b9ddb8a6311bff6f5e29cb3722d1f4236d66292
//Author: Haoyuan Feng <fenghaoyuan19@mails.ucas.ac.cn>
//Date:   Mon Feb 10 11:08:16 2025 +0800
//
//    fix(MMU): Should consider s2xlate when calculate page level (#4253)
//diff --git a/.gitignore b/.gitignore
//index 09907c997..39a1a9ef4 100644
//--- a/.gitignore
//+++ b/.gitignore
//@@ -288,7 +288,6 @@ Temporary Items
// # gitignore contributors: remember to update Global/Xcode.gitignore, Objective-C.gitignore & Swift.gitignore
// 
// ## Build generated
//-build
// DerivedData
// 
// ## Various settings
// Generated by CIRCT firtool-1.62.1
// Standard header to adapt well known macros for register randomization.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module XSTop(
  input          nmi_0_0,
  input          nmi_0_1,
  output         dma_awready,
  input          dma_awvalid,
  input  [13:0]  dma_awid,
  input  [47:0]  dma_awaddr,
  input  [7:0]   dma_awlen,
  input  [2:0]   dma_awsize,
  input  [1:0]   dma_awburst,
  input          dma_awlock,
  input  [3:0]   dma_awcache,
  input  [2:0]   dma_awprot,
  input  [3:0]   dma_awqos,
  output         dma_wready,
  input          dma_wvalid,
  input  [255:0] dma_wdata,
  input  [31:0]  dma_wstrb,
  input          dma_wlast,
  input          dma_bready,
  output         dma_bvalid,
  output [13:0]  dma_bid,
  output [1:0]   dma_bresp,
  output         dma_arready,
  input          dma_arvalid,
  input  [13:0]  dma_arid,
  input  [47:0]  dma_araddr,
  input  [7:0]   dma_arlen,
  input  [2:0]   dma_arsize,
  input  [1:0]   dma_arburst,
  input          dma_arlock,
  input  [3:0]   dma_arcache,
  input  [2:0]   dma_arprot,
  input  [3:0]   dma_arqos,
  input          dma_rready,
  output         dma_rvalid,
  output [13:0]  dma_rid,
  output [255:0] dma_rdata,
  output [1:0]   dma_rresp,
  output         dma_rlast,
  input          peripheral_awready,
  output         peripheral_awvalid,
  output [1:0]   peripheral_awid,
  output [30:0]  peripheral_awaddr,
  output [7:0]   peripheral_awlen,
  output [2:0]   peripheral_awsize,
  output [1:0]   peripheral_awburst,
  output         peripheral_awlock,
  output [3:0]   peripheral_awcache,
  output [2:0]   peripheral_awprot,
  output [3:0]   peripheral_awqos,
  input          peripheral_wready,
  output         peripheral_wvalid,
  output [63:0]  peripheral_wdata,
  output [7:0]   peripheral_wstrb,
  output         peripheral_wlast,
  output         peripheral_bready,
  input          peripheral_bvalid,
  input  [1:0]   peripheral_bid,
  input  [1:0]   peripheral_bresp,
  input          peripheral_arready,
  output         peripheral_arvalid,
  output [1:0]   peripheral_arid,
  output [30:0]  peripheral_araddr,
  output [7:0]   peripheral_arlen,
  output [2:0]   peripheral_arsize,
  output [1:0]   peripheral_arburst,
  output         peripheral_arlock,
  output [3:0]   peripheral_arcache,
  output [2:0]   peripheral_arprot,
  output [3:0]   peripheral_arqos,
  output         peripheral_rready,
  input          peripheral_rvalid,
  input  [1:0]   peripheral_rid,
  input  [63:0]  peripheral_rdata,
  input  [1:0]   peripheral_rresp,
  input          peripheral_rlast,
  input          memory_awready,
  output         memory_awvalid,
  output [13:0]  memory_awid,
  output [47:0]  memory_awaddr,
  output [7:0]   memory_awlen,
  output [2:0]   memory_awsize,
  output [1:0]   memory_awburst,
  output         memory_awlock,
  output [3:0]   memory_awcache,
  output [2:0]   memory_awprot,
  output [3:0]   memory_awqos,
  input          memory_wready,
  output         memory_wvalid,
  output [255:0] memory_wdata,
  output [31:0]  memory_wstrb,
  output         memory_wlast,
  output         memory_bready,
  input          memory_bvalid,
  input  [13:0]  memory_bid,
  input  [1:0]   memory_bresp,
  input          memory_arready,
  output         memory_arvalid,
  output [13:0]  memory_arid,
  output [47:0]  memory_araddr,
  output [7:0]   memory_arlen,
  output [2:0]   memory_arsize,
  output [1:0]   memory_arburst,
  output         memory_arlock,
  output [3:0]   memory_arcache,
  output [2:0]   memory_arprot,
  output [3:0]   memory_arqos,
  output         memory_rready,
  input          memory_rvalid,
  input  [13:0]  memory_rid,
  input  [255:0] memory_rdata,
  input  [1:0]   memory_rresp,
  input          memory_rlast,
  input          io_clock,
  input          io_reset,
  input  [15:0]  io_sram_config,
  input  [63:0]  io_extIntrs,
  input          io_pll0_lock,
  output [31:0]  io_pll0_ctrl_0,
  output [31:0]  io_pll0_ctrl_1,
  output [31:0]  io_pll0_ctrl_2,
  output [31:0]  io_pll0_ctrl_3,
  output [31:0]  io_pll0_ctrl_4,
  output [31:0]  io_pll0_ctrl_5,
  input          io_systemjtag_jtag_TCK,
  input          io_systemjtag_jtag_TMS,
  input          io_systemjtag_jtag_TDI,
  output         io_systemjtag_jtag_TDO_data,
  output         io_systemjtag_jtag_TDO_driven,
  input          io_systemjtag_reset,
  input  [10:0]  io_systemjtag_mfr_id,
  input  [15:0]  io_systemjtag_part_number,
  input  [3:0]   io_systemjtag_version,
  output         io_debug_reset,
  input          io_rtc_clock,
  input          io_cacheable_check_req_0_valid,
  input  [47:0]  io_cacheable_check_req_0_bits_addr,
  input  [1:0]   io_cacheable_check_req_0_bits_size,
  input  [2:0]   io_cacheable_check_req_0_bits_cmd,
  input          io_cacheable_check_req_1_valid,
  input  [47:0]  io_cacheable_check_req_1_bits_addr,
  input  [1:0]   io_cacheable_check_req_1_bits_size,
  input  [2:0]   io_cacheable_check_req_1_bits_cmd,
  output         io_cacheable_check_resp_0_ld,
  output         io_cacheable_check_resp_0_st,
  output         io_cacheable_check_resp_0_instr,
  output         io_cacheable_check_resp_0_mmio,
  output         io_cacheable_check_resp_0_atomic,
  output         io_cacheable_check_resp_1_ld,
  output         io_cacheable_check_resp_1_st,
  output         io_cacheable_check_resp_1_instr,
  output         io_cacheable_check_resp_1_mmio,
  output         io_cacheable_check_resp_1_atomic,
  output         io_riscv_halt_0,
  output         io_riscv_critical_error_0,
  input  [47:0]  io_riscv_rst_vec_0,
  input          io_traceCoreInterface_0_fromEncoder_enable,
  input          io_traceCoreInterface_0_fromEncoder_stall,
  output [63:0]  io_traceCoreInterface_0_toEncoder_cause,
  output [49:0]  io_traceCoreInterface_0_toEncoder_tval,
  output [2:0]   io_traceCoreInterface_0_toEncoder_priv,
  output [149:0] io_traceCoreInterface_0_toEncoder_iaddr,
  output [11:0]  io_traceCoreInterface_0_toEncoder_itype,
  output [20:0]  io_traceCoreInterface_0_toEncoder_iretire,
  output [2:0]   io_traceCoreInterface_0_toEncoder_ilastsize
);

  wire         _resetGen_1_o_reset;
  wire         _resetGen_o_reset;
  wire         _jtag_reset_sync_resetSync_o_reset;
  wire         _reset_sync_resetSync_o_reset;
  wire         _broadcast_auto_out_valid;
  wire [5:0]   _broadcast_auto_out_bits_hartid;
  wire [41:0]  _broadcast_auto_out_bits_rawData_0;
  wire [41:0]  _broadcast_auto_out_bits_rawData_1;
  wire [41:0]  _broadcast_auto_out_bits_rawData_2;
  wire         _intBuffer_1_auto_out_0;
  wire         _intBuffer_auto_out_0;
  wire         _l3cacheOpt_auto_ctrl_unit_int_out_0;
  wire         _l3cacheOpt_auto_ctrl_unit_ctl_in_a_ready;
  wire         _l3cacheOpt_auto_ctrl_unit_ctl_in_d_valid;
  wire [3:0]   _l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_opcode;
  wire [1:0]   _l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_size;
  wire [2:0]   _l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_source;
  wire [63:0]  _l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_data;
  wire         _l3cacheOpt_auto_tpmeta_send_out_valid;
  wire [5:0]   _l3cacheOpt_auto_tpmeta_send_out_bits_hartid;
  wire [41:0]  _l3cacheOpt_auto_tpmeta_send_out_bits_rawData_0;
  wire [41:0]  _l3cacheOpt_auto_tpmeta_send_out_bits_rawData_1;
  wire [41:0]  _l3cacheOpt_auto_tpmeta_send_out_bits_rawData_2;
  wire         _l3cacheOpt_auto_tpmeta_recv_in_ready;
  wire         _l3cacheOpt_auto_in_a_ready;
  wire         _l3cacheOpt_auto_in_b_valid;
  wire [1:0]   _l3cacheOpt_auto_in_b_bits_param;
  wire [47:0]  _l3cacheOpt_auto_in_b_bits_address;
  wire [255:0] _l3cacheOpt_auto_in_b_bits_data;
  wire         _l3cacheOpt_auto_in_c_ready;
  wire         _l3cacheOpt_auto_in_d_valid;
  wire [3:0]   _l3cacheOpt_auto_in_d_bits_opcode;
  wire [1:0]   _l3cacheOpt_auto_in_d_bits_param;
  wire [2:0]   _l3cacheOpt_auto_in_d_bits_size;
  wire [10:0]  _l3cacheOpt_auto_in_d_bits_source;
  wire [3:0]   _l3cacheOpt_auto_in_d_bits_sink;
  wire         _l3cacheOpt_auto_in_d_bits_denied;
  wire         _l3cacheOpt_auto_in_d_bits_echo_blockisdirty;
  wire [255:0] _l3cacheOpt_auto_in_d_bits_data;
  wire         _l3cacheOpt_auto_in_d_bits_corrupt;
  wire         _l3cacheOpt_auto_out_a_valid;
  wire [3:0]   _l3cacheOpt_auto_out_a_bits_opcode;
  wire [2:0]   _l3cacheOpt_auto_out_a_bits_param;
  wire [2:0]   _l3cacheOpt_auto_out_a_bits_size;
  wire [3:0]   _l3cacheOpt_auto_out_a_bits_source;
  wire [47:0]  _l3cacheOpt_auto_out_a_bits_address;
  wire [31:0]  _l3cacheOpt_auto_out_a_bits_mask;
  wire [255:0] _l3cacheOpt_auto_out_a_bits_data;
  wire         _l3cacheOpt_auto_out_a_bits_corrupt;
  wire         _l3cacheOpt_auto_out_c_valid;
  wire [2:0]   _l3cacheOpt_auto_out_c_bits_opcode;
  wire [2:0]   _l3cacheOpt_auto_out_c_bits_size;
  wire [3:0]   _l3cacheOpt_auto_out_c_bits_source;
  wire [47:0]  _l3cacheOpt_auto_out_c_bits_address;
  wire [255:0] _l3cacheOpt_auto_out_c_bits_data;
  wire         _l3cacheOpt_auto_out_c_bits_corrupt;
  wire         _l3cacheOpt_auto_out_d_ready;
  wire         _l3cacheOpt_auto_out_e_valid;
  wire [2:0]   _l3cacheOpt_auto_out_e_bits_sink;
  wire         _l3cacheOpt_io_l3Miss;
  wire         _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_valid;
  wire [5:0]   _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_hartid;
  wire [31:0]  _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_set;
  wire [3:0]   _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_way;
  wire         _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_wmode;
  wire [41:0]  _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_0;
  wire [41:0]  _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_1;
  wire [41:0]  _core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_2;
  wire         _core_with_l2_auto_l2top_inner_beu_int_out_0;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_a_valid;
  wire [3:0]   _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_opcode;
  wire [2:0]   _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_param;
  wire [2:0]   _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_size;
  wire [9:0]   _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_source;
  wire [47:0]  _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_address;
  wire [3:0]   _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_user_reqSource;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_echo_blockisdirty;
  wire [31:0]  _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_mask;
  wire [255:0] _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_data;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_a_bits_corrupt;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_b_ready;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_c_valid;
  wire [2:0]   _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_opcode;
  wire [2:0]   _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_param;
  wire [2:0]   _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_size;
  wire [9:0]   _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_source;
  wire [47:0]  _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_address;
  wire [3:0]   _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_user_reqSource;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_echo_blockisdirty;
  wire [255:0] _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_data;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_c_bits_corrupt;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_d_ready;
  wire         _core_with_l2_auto_l2top_inner_memory_port_out_e_valid;
  wire [3:0]   _core_with_l2_auto_l2top_inner_memory_port_out_e_bits_sink;
  wire         _core_with_l2_auto_l2top_inner_mmio_port_out_a_valid;
  wire [3:0]   _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_opcode;
  wire [2:0]   _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_param;
  wire [2:0]   _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_size;
  wire [2:0]   _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_source;
  wire [47:0]  _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_address;
  wire [7:0]   _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_mask;
  wire [63:0]  _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_data;
  wire         _core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_corrupt;
  wire         _core_with_l2_auto_l2top_inner_mmio_port_out_d_ready;
  wire [63:0]  _core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr;
  wire         _core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr_valid;
  wire         _core_with_l2_io_hartIsInReset;
  wire [49:0]  _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iaddr;
  wire [3:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_itype;
  wire [6:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iretire;
  wire         _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_ilastsize;
  wire [49:0]  _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iaddr;
  wire [3:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_itype;
  wire [6:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iretire;
  wire         _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_ilastsize;
  wire [49:0]  _core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iaddr;
  wire [3:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_itype;
  wire [6:0]   _core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iretire;
  wire         _core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_ilastsize;
  wire         _socMisc_auto_debugModule_debug_dmOuter_dmOuter_int_out_0;
  wire         _socMisc_auto_plic_int_out_1_0;
  wire         _socMisc_auto_plic_int_out_0_0;
  wire         _socMisc_auto_clint_int_out_0;
  wire         _socMisc_auto_clint_int_out_1;
  wire         _socMisc_auto_buffer_in_a_ready;
  wire         _socMisc_auto_buffer_in_b_valid;
  wire [2:0]   _socMisc_auto_buffer_in_b_bits_opcode;
  wire [1:0]   _socMisc_auto_buffer_in_b_bits_param;
  wire [2:0]   _socMisc_auto_buffer_in_b_bits_size;
  wire [47:0]  _socMisc_auto_buffer_in_b_bits_address;
  wire [31:0]  _socMisc_auto_buffer_in_b_bits_mask;
  wire [255:0] _socMisc_auto_buffer_in_b_bits_data;
  wire         _socMisc_auto_buffer_in_b_bits_corrupt;
  wire         _socMisc_auto_buffer_in_c_ready;
  wire         _socMisc_auto_buffer_in_d_valid;
  wire [3:0]   _socMisc_auto_buffer_in_d_bits_opcode;
  wire [1:0]   _socMisc_auto_buffer_in_d_bits_param;
  wire [2:0]   _socMisc_auto_buffer_in_d_bits_size;
  wire [9:0]   _socMisc_auto_buffer_in_d_bits_source;
  wire [3:0]   _socMisc_auto_buffer_in_d_bits_sink;
  wire         _socMisc_auto_buffer_in_d_bits_denied;
  wire         _socMisc_auto_buffer_in_d_bits_echo_blockisdirty;
  wire [255:0] _socMisc_auto_buffer_in_d_bits_data;
  wire         _socMisc_auto_buffer_in_d_bits_corrupt;
  wire         _socMisc_auto_buffer_in_e_ready;
  wire         _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_a_ready;
  wire         _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_valid;
  wire [3:0]   _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_opcode;
  wire [1:0]   _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_param;
  wire [2:0]   _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_size;
  wire [2:0]   _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_source;
  wire         _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_sink;
  wire         _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_denied;
  wire [63:0]  _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_data;
  wire         _socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_corrupt;
  wire         _socMisc_auto_xbar_out_1_a_valid;
  wire [3:0]   _socMisc_auto_xbar_out_1_a_bits_opcode;
  wire [2:0]   _socMisc_auto_xbar_out_1_a_bits_param;
  wire [2:0]   _socMisc_auto_xbar_out_1_a_bits_size;
  wire [10:0]  _socMisc_auto_xbar_out_1_a_bits_source;
  wire [47:0]  _socMisc_auto_xbar_out_1_a_bits_address;
  wire [3:0]   _socMisc_auto_xbar_out_1_a_bits_user_reqSource;
  wire [31:0]  _socMisc_auto_xbar_out_1_a_bits_mask;
  wire [255:0] _socMisc_auto_xbar_out_1_a_bits_data;
  wire         _socMisc_auto_xbar_out_1_a_bits_corrupt;
  wire         _socMisc_auto_xbar_out_1_b_ready;
  wire         _socMisc_auto_xbar_out_1_c_valid;
  wire [2:0]   _socMisc_auto_xbar_out_1_c_bits_opcode;
  wire [2:0]   _socMisc_auto_xbar_out_1_c_bits_param;
  wire [2:0]   _socMisc_auto_xbar_out_1_c_bits_size;
  wire [10:0]  _socMisc_auto_xbar_out_1_c_bits_source;
  wire [47:0]  _socMisc_auto_xbar_out_1_c_bits_address;
  wire         _socMisc_auto_xbar_out_1_c_bits_echo_blockisdirty;
  wire [255:0] _socMisc_auto_xbar_out_1_c_bits_data;
  wire         _socMisc_auto_xbar_out_1_d_ready;
  wire         _socMisc_auto_xbar_out_1_e_valid;
  wire [3:0]   _socMisc_auto_xbar_out_1_e_bits_sink;
  wire         _socMisc_auto_xbar_out_0_a_valid;
  wire [3:0]   _socMisc_auto_xbar_out_0_a_bits_opcode;
  wire [1:0]   _socMisc_auto_xbar_out_0_a_bits_size;
  wire [2:0]   _socMisc_auto_xbar_out_0_a_bits_source;
  wire [29:0]  _socMisc_auto_xbar_out_0_a_bits_address;
  wire [7:0]   _socMisc_auto_xbar_out_0_a_bits_mask;
  wire [63:0]  _socMisc_auto_xbar_out_0_a_bits_data;
  wire         _socMisc_auto_xbar_out_0_d_ready;
  wire         _socMisc_auto_binder_in_a_ready;
  wire         _socMisc_auto_binder_in_c_ready;
  wire         _socMisc_auto_binder_in_d_valid;
  wire [3:0]   _socMisc_auto_binder_in_d_bits_opcode;
  wire [1:0]   _socMisc_auto_binder_in_d_bits_param;
  wire [2:0]   _socMisc_auto_binder_in_d_bits_size;
  wire [3:0]   _socMisc_auto_binder_in_d_bits_source;
  wire [2:0]   _socMisc_auto_binder_in_d_bits_sink;
  wire         _socMisc_auto_binder_in_d_bits_denied;
  wire [255:0] _socMisc_auto_binder_in_d_bits_data;
  wire         _socMisc_auto_binder_in_d_bits_corrupt;
  wire         _socMisc_debug_module_io_resetCtrl_hartResetReq_0;
  wire         _socMisc_debug_module_io_debugIO_dmactive;
  wire         _socMisc_clintTime_valid;
  wire [63:0]  _socMisc_clintTime_bits;
  SoCMisc socMisc (
    .clock                                               (io_clock),
    .reset                                               (_resetGen_o_reset),
    .auto_debugModule_debug_dmOuter_dmOuter_int_out_0
      (_socMisc_auto_debugModule_debug_dmOuter_dmOuter_int_out_0),
    .auto_plic_int_in_1_0                                (_intBuffer_1_auto_out_0),
    .auto_plic_int_in_0_0                                (_intBuffer_auto_out_0),
    .auto_plic_int_out_1_0                               (_socMisc_auto_plic_int_out_1_0),
    .auto_plic_int_out_0_0                               (_socMisc_auto_plic_int_out_0_0),
    .auto_clint_int_out_0                                (_socMisc_auto_clint_int_out_0),
    .auto_clint_int_out_1                                (_socMisc_auto_clint_int_out_1),
    .auto_buffer_in_a_ready
      (_socMisc_auto_buffer_in_a_ready),
    .auto_buffer_in_a_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_valid),
    .auto_buffer_in_a_bits_opcode
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_opcode),
    .auto_buffer_in_a_bits_param
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_param),
    .auto_buffer_in_a_bits_size
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_size),
    .auto_buffer_in_a_bits_source
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_source),
    .auto_buffer_in_a_bits_address
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_address),
    .auto_buffer_in_a_bits_user_reqSource
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_user_reqSource),
    .auto_buffer_in_a_bits_echo_blockisdirty
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_echo_blockisdirty),
    .auto_buffer_in_a_bits_mask
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_mask),
    .auto_buffer_in_a_bits_data
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_data),
    .auto_buffer_in_a_bits_corrupt
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_corrupt),
    .auto_buffer_in_b_ready
      (_core_with_l2_auto_l2top_inner_memory_port_out_b_ready),
    .auto_buffer_in_b_valid
      (_socMisc_auto_buffer_in_b_valid),
    .auto_buffer_in_b_bits_opcode
      (_socMisc_auto_buffer_in_b_bits_opcode),
    .auto_buffer_in_b_bits_param
      (_socMisc_auto_buffer_in_b_bits_param),
    .auto_buffer_in_b_bits_size
      (_socMisc_auto_buffer_in_b_bits_size),
    .auto_buffer_in_b_bits_address
      (_socMisc_auto_buffer_in_b_bits_address),
    .auto_buffer_in_b_bits_mask
      (_socMisc_auto_buffer_in_b_bits_mask),
    .auto_buffer_in_b_bits_data
      (_socMisc_auto_buffer_in_b_bits_data),
    .auto_buffer_in_b_bits_corrupt
      (_socMisc_auto_buffer_in_b_bits_corrupt),
    .auto_buffer_in_c_ready
      (_socMisc_auto_buffer_in_c_ready),
    .auto_buffer_in_c_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_valid),
    .auto_buffer_in_c_bits_opcode
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_opcode),
    .auto_buffer_in_c_bits_param
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_param),
    .auto_buffer_in_c_bits_size
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_size),
    .auto_buffer_in_c_bits_source
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_source),
    .auto_buffer_in_c_bits_address
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_address),
    .auto_buffer_in_c_bits_user_reqSource
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_user_reqSource),
    .auto_buffer_in_c_bits_echo_blockisdirty
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_echo_blockisdirty),
    .auto_buffer_in_c_bits_data
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_data),
    .auto_buffer_in_c_bits_corrupt
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_corrupt),
    .auto_buffer_in_d_ready
      (_core_with_l2_auto_l2top_inner_memory_port_out_d_ready),
    .auto_buffer_in_d_valid
      (_socMisc_auto_buffer_in_d_valid),
    .auto_buffer_in_d_bits_opcode
      (_socMisc_auto_buffer_in_d_bits_opcode),
    .auto_buffer_in_d_bits_param
      (_socMisc_auto_buffer_in_d_bits_param),
    .auto_buffer_in_d_bits_size
      (_socMisc_auto_buffer_in_d_bits_size),
    .auto_buffer_in_d_bits_source
      (_socMisc_auto_buffer_in_d_bits_source),
    .auto_buffer_in_d_bits_sink
      (_socMisc_auto_buffer_in_d_bits_sink),
    .auto_buffer_in_d_bits_denied
      (_socMisc_auto_buffer_in_d_bits_denied),
    .auto_buffer_in_d_bits_echo_blockisdirty
      (_socMisc_auto_buffer_in_d_bits_echo_blockisdirty),
    .auto_buffer_in_d_bits_data
      (_socMisc_auto_buffer_in_d_bits_data),
    .auto_buffer_in_d_bits_corrupt
      (_socMisc_auto_buffer_in_d_bits_corrupt),
    .auto_buffer_in_e_ready
      (_socMisc_auto_buffer_in_e_ready),
    .auto_buffer_in_e_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_e_valid),
    .auto_buffer_in_e_bits_sink
      (_core_with_l2_auto_l2top_inner_memory_port_out_e_bits_sink),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_ready
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_a_ready),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_valid
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_valid),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_opcode
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_opcode),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_param
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_param),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_size
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_size),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_source
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_source),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_address
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_address),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_mask
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_mask),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_data
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_data),
    .auto_L2_to_L3_peripheral_buffer_1_in_a_bits_corrupt
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_corrupt),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_ready
      (_core_with_l2_auto_l2top_inner_mmio_port_out_d_ready),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_valid
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_valid),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_opcode
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_opcode),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_param
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_param),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_size
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_size),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_source
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_source),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_sink
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_sink),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_denied
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_denied),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_data
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_data),
    .auto_L2_to_L3_peripheral_buffer_1_in_d_bits_corrupt
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_corrupt),
    .auto_xbar_out_1_a_ready                             (_l3cacheOpt_auto_in_a_ready),
    .auto_xbar_out_1_a_valid
      (_socMisc_auto_xbar_out_1_a_valid),
    .auto_xbar_out_1_a_bits_opcode
      (_socMisc_auto_xbar_out_1_a_bits_opcode),
    .auto_xbar_out_1_a_bits_param
      (_socMisc_auto_xbar_out_1_a_bits_param),
    .auto_xbar_out_1_a_bits_size
      (_socMisc_auto_xbar_out_1_a_bits_size),
    .auto_xbar_out_1_a_bits_source
      (_socMisc_auto_xbar_out_1_a_bits_source),
    .auto_xbar_out_1_a_bits_address
      (_socMisc_auto_xbar_out_1_a_bits_address),
    .auto_xbar_out_1_a_bits_user_reqSource
      (_socMisc_auto_xbar_out_1_a_bits_user_reqSource),
    .auto_xbar_out_1_a_bits_mask
      (_socMisc_auto_xbar_out_1_a_bits_mask),
    .auto_xbar_out_1_a_bits_data
      (_socMisc_auto_xbar_out_1_a_bits_data),
    .auto_xbar_out_1_a_bits_corrupt
      (_socMisc_auto_xbar_out_1_a_bits_corrupt),
    .auto_xbar_out_1_b_ready
      (_socMisc_auto_xbar_out_1_b_ready),
    .auto_xbar_out_1_b_valid                             (_l3cacheOpt_auto_in_b_valid),
    .auto_xbar_out_1_b_bits_param
      (_l3cacheOpt_auto_in_b_bits_param),
    .auto_xbar_out_1_b_bits_address
      (_l3cacheOpt_auto_in_b_bits_address),
    .auto_xbar_out_1_b_bits_data
      (_l3cacheOpt_auto_in_b_bits_data),
    .auto_xbar_out_1_c_ready                             (_l3cacheOpt_auto_in_c_ready),
    .auto_xbar_out_1_c_valid
      (_socMisc_auto_xbar_out_1_c_valid),
    .auto_xbar_out_1_c_bits_opcode
      (_socMisc_auto_xbar_out_1_c_bits_opcode),
    .auto_xbar_out_1_c_bits_param
      (_socMisc_auto_xbar_out_1_c_bits_param),
    .auto_xbar_out_1_c_bits_size
      (_socMisc_auto_xbar_out_1_c_bits_size),
    .auto_xbar_out_1_c_bits_source
      (_socMisc_auto_xbar_out_1_c_bits_source),
    .auto_xbar_out_1_c_bits_address
      (_socMisc_auto_xbar_out_1_c_bits_address),
    .auto_xbar_out_1_c_bits_echo_blockisdirty
      (_socMisc_auto_xbar_out_1_c_bits_echo_blockisdirty),
    .auto_xbar_out_1_c_bits_data
      (_socMisc_auto_xbar_out_1_c_bits_data),
    .auto_xbar_out_1_d_ready
      (_socMisc_auto_xbar_out_1_d_ready),
    .auto_xbar_out_1_d_valid                             (_l3cacheOpt_auto_in_d_valid),
    .auto_xbar_out_1_d_bits_opcode
      (_l3cacheOpt_auto_in_d_bits_opcode),
    .auto_xbar_out_1_d_bits_param
      (_l3cacheOpt_auto_in_d_bits_param),
    .auto_xbar_out_1_d_bits_size
      (_l3cacheOpt_auto_in_d_bits_size),
    .auto_xbar_out_1_d_bits_source
      (_l3cacheOpt_auto_in_d_bits_source),
    .auto_xbar_out_1_d_bits_sink
      (_l3cacheOpt_auto_in_d_bits_sink),
    .auto_xbar_out_1_d_bits_denied
      (_l3cacheOpt_auto_in_d_bits_denied),
    .auto_xbar_out_1_d_bits_echo_blockisdirty
      (_l3cacheOpt_auto_in_d_bits_echo_blockisdirty),
    .auto_xbar_out_1_d_bits_data
      (_l3cacheOpt_auto_in_d_bits_data),
    .auto_xbar_out_1_d_bits_corrupt
      (_l3cacheOpt_auto_in_d_bits_corrupt),
    .auto_xbar_out_1_e_valid
      (_socMisc_auto_xbar_out_1_e_valid),
    .auto_xbar_out_1_e_bits_sink
      (_socMisc_auto_xbar_out_1_e_bits_sink),
    .auto_xbar_out_0_a_ready
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_a_ready),
    .auto_xbar_out_0_a_valid
      (_socMisc_auto_xbar_out_0_a_valid),
    .auto_xbar_out_0_a_bits_opcode
      (_socMisc_auto_xbar_out_0_a_bits_opcode),
    .auto_xbar_out_0_a_bits_size
      (_socMisc_auto_xbar_out_0_a_bits_size),
    .auto_xbar_out_0_a_bits_source
      (_socMisc_auto_xbar_out_0_a_bits_source),
    .auto_xbar_out_0_a_bits_address
      (_socMisc_auto_xbar_out_0_a_bits_address),
    .auto_xbar_out_0_a_bits_mask
      (_socMisc_auto_xbar_out_0_a_bits_mask),
    .auto_xbar_out_0_a_bits_data
      (_socMisc_auto_xbar_out_0_a_bits_data),
    .auto_xbar_out_0_d_ready
      (_socMisc_auto_xbar_out_0_d_ready),
    .auto_xbar_out_0_d_valid
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_valid),
    .auto_xbar_out_0_d_bits_opcode
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_opcode),
    .auto_xbar_out_0_d_bits_size
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_size),
    .auto_xbar_out_0_d_bits_source
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_source),
    .auto_xbar_out_0_d_bits_data
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_data),
    .auto_binder_in_a_ready
      (_socMisc_auto_binder_in_a_ready),
    .auto_binder_in_a_valid                              (_l3cacheOpt_auto_out_a_valid),
    .auto_binder_in_a_bits_opcode
      (_l3cacheOpt_auto_out_a_bits_opcode),
    .auto_binder_in_a_bits_param
      (_l3cacheOpt_auto_out_a_bits_param),
    .auto_binder_in_a_bits_size
      (_l3cacheOpt_auto_out_a_bits_size),
    .auto_binder_in_a_bits_source
      (_l3cacheOpt_auto_out_a_bits_source),
    .auto_binder_in_a_bits_address
      (_l3cacheOpt_auto_out_a_bits_address),
    .auto_binder_in_a_bits_mask
      (_l3cacheOpt_auto_out_a_bits_mask),
    .auto_binder_in_a_bits_data
      (_l3cacheOpt_auto_out_a_bits_data),
    .auto_binder_in_a_bits_corrupt
      (_l3cacheOpt_auto_out_a_bits_corrupt),
    .auto_binder_in_c_ready
      (_socMisc_auto_binder_in_c_ready),
    .auto_binder_in_c_valid                              (_l3cacheOpt_auto_out_c_valid),
    .auto_binder_in_c_bits_opcode
      (_l3cacheOpt_auto_out_c_bits_opcode),
    .auto_binder_in_c_bits_size
      (_l3cacheOpt_auto_out_c_bits_size),
    .auto_binder_in_c_bits_source
      (_l3cacheOpt_auto_out_c_bits_source),
    .auto_binder_in_c_bits_address
      (_l3cacheOpt_auto_out_c_bits_address),
    .auto_binder_in_c_bits_data
      (_l3cacheOpt_auto_out_c_bits_data),
    .auto_binder_in_c_bits_corrupt
      (_l3cacheOpt_auto_out_c_bits_corrupt),
    .auto_binder_in_d_ready                              (_l3cacheOpt_auto_out_d_ready),
    .auto_binder_in_d_valid
      (_socMisc_auto_binder_in_d_valid),
    .auto_binder_in_d_bits_opcode
      (_socMisc_auto_binder_in_d_bits_opcode),
    .auto_binder_in_d_bits_param
      (_socMisc_auto_binder_in_d_bits_param),
    .auto_binder_in_d_bits_size
      (_socMisc_auto_binder_in_d_bits_size),
    .auto_binder_in_d_bits_source
      (_socMisc_auto_binder_in_d_bits_source),
    .auto_binder_in_d_bits_sink
      (_socMisc_auto_binder_in_d_bits_sink),
    .auto_binder_in_d_bits_denied
      (_socMisc_auto_binder_in_d_bits_denied),
    .auto_binder_in_d_bits_data
      (_socMisc_auto_binder_in_d_bits_data),
    .auto_binder_in_d_bits_corrupt
      (_socMisc_auto_binder_in_d_bits_corrupt),
    .auto_binder_in_e_valid                              (_l3cacheOpt_auto_out_e_valid),
    .auto_binder_in_e_bits_sink
      (_l3cacheOpt_auto_out_e_bits_sink),
    .memory_0_aw_ready                                   (memory_awready),
    .memory_0_aw_valid                                   (memory_awvalid),
    .memory_0_aw_bits_id                                 (memory_awid),
    .memory_0_aw_bits_addr                               (memory_awaddr),
    .memory_0_aw_bits_len                                (memory_awlen),
    .memory_0_aw_bits_size                               (memory_awsize),
    .memory_0_aw_bits_burst                              (memory_awburst),
    .memory_0_aw_bits_lock                               (memory_awlock),
    .memory_0_aw_bits_cache                              (memory_awcache),
    .memory_0_aw_bits_prot                               (memory_awprot),
    .memory_0_aw_bits_qos                                (memory_awqos),
    .memory_0_w_ready                                    (memory_wready),
    .memory_0_w_valid                                    (memory_wvalid),
    .memory_0_w_bits_data                                (memory_wdata),
    .memory_0_w_bits_strb                                (memory_wstrb),
    .memory_0_w_bits_last                                (memory_wlast),
    .memory_0_b_ready                                    (memory_bready),
    .memory_0_b_valid                                    (memory_bvalid),
    .memory_0_b_bits_id                                  (memory_bid),
    .memory_0_b_bits_resp                                (memory_bresp),
    .memory_0_ar_ready                                   (memory_arready),
    .memory_0_ar_valid                                   (memory_arvalid),
    .memory_0_ar_bits_id                                 (memory_arid),
    .memory_0_ar_bits_addr                               (memory_araddr),
    .memory_0_ar_bits_len                                (memory_arlen),
    .memory_0_ar_bits_size                               (memory_arsize),
    .memory_0_ar_bits_burst                              (memory_arburst),
    .memory_0_ar_bits_lock                               (memory_arlock),
    .memory_0_ar_bits_cache                              (memory_arcache),
    .memory_0_ar_bits_prot                               (memory_arprot),
    .memory_0_ar_bits_qos                                (memory_arqos),
    .memory_0_r_ready                                    (memory_rready),
    .memory_0_r_valid                                    (memory_rvalid),
    .memory_0_r_bits_id                                  (memory_rid),
    .memory_0_r_bits_data                                (memory_rdata),
    .memory_0_r_bits_resp                                (memory_rresp),
    .memory_0_r_bits_last                                (memory_rlast),
    .peripheral_0_aw_ready                               (peripheral_awready),
    .peripheral_0_aw_valid                               (peripheral_awvalid),
    .peripheral_0_aw_bits_id                             (peripheral_awid),
    .peripheral_0_aw_bits_addr                           (peripheral_awaddr),
    .peripheral_0_aw_bits_len                            (peripheral_awlen),
    .peripheral_0_aw_bits_size                           (peripheral_awsize),
    .peripheral_0_aw_bits_burst                          (peripheral_awburst),
    .peripheral_0_aw_bits_lock                           (peripheral_awlock),
    .peripheral_0_aw_bits_cache                          (peripheral_awcache),
    .peripheral_0_aw_bits_prot                           (peripheral_awprot),
    .peripheral_0_aw_bits_qos                            (peripheral_awqos),
    .peripheral_0_w_ready                                (peripheral_wready),
    .peripheral_0_w_valid                                (peripheral_wvalid),
    .peripheral_0_w_bits_data                            (peripheral_wdata),
    .peripheral_0_w_bits_strb                            (peripheral_wstrb),
    .peripheral_0_w_bits_last                            (peripheral_wlast),
    .peripheral_0_b_ready                                (peripheral_bready),
    .peripheral_0_b_valid                                (peripheral_bvalid),
    .peripheral_0_b_bits_id                              (peripheral_bid),
    .peripheral_0_b_bits_resp                            (peripheral_bresp),
    .peripheral_0_ar_ready                               (peripheral_arready),
    .peripheral_0_ar_valid                               (peripheral_arvalid),
    .peripheral_0_ar_bits_id                             (peripheral_arid),
    .peripheral_0_ar_bits_addr                           (peripheral_araddr),
    .peripheral_0_ar_bits_len                            (peripheral_arlen),
    .peripheral_0_ar_bits_size                           (peripheral_arsize),
    .peripheral_0_ar_bits_burst                          (peripheral_arburst),
    .peripheral_0_ar_bits_lock                           (peripheral_arlock),
    .peripheral_0_ar_bits_cache                          (peripheral_arcache),
    .peripheral_0_ar_bits_prot                           (peripheral_arprot),
    .peripheral_0_ar_bits_qos                            (peripheral_arqos),
    .peripheral_0_r_ready                                (peripheral_rready),
    .peripheral_0_r_valid                                (peripheral_rvalid),
    .peripheral_0_r_bits_id                              (peripheral_rid),
    .peripheral_0_r_bits_data                            (peripheral_rdata),
    .peripheral_0_r_bits_resp                            (peripheral_rresp),
    .peripheral_0_r_bits_last                            (peripheral_rlast),
    .dma_0_aw_ready                                      (dma_awready),
    .dma_0_aw_valid                                      (dma_awvalid),
    .dma_0_aw_bits_id                                    (dma_awid),
    .dma_0_aw_bits_addr                                  (dma_awaddr),
    .dma_0_aw_bits_len                                   (dma_awlen),
    .dma_0_aw_bits_size                                  (dma_awsize),
    .dma_0_aw_bits_burst                                 (dma_awburst),
    .dma_0_aw_bits_lock                                  (dma_awlock),
    .dma_0_aw_bits_cache                                 (dma_awcache),
    .dma_0_aw_bits_prot                                  (dma_awprot),
    .dma_0_aw_bits_qos                                   (dma_awqos),
    .dma_0_w_ready                                       (dma_wready),
    .dma_0_w_valid                                       (dma_wvalid),
    .dma_0_w_bits_data                                   (dma_wdata),
    .dma_0_w_bits_strb                                   (dma_wstrb),
    .dma_0_w_bits_last                                   (dma_wlast),
    .dma_0_b_ready                                       (dma_bready),
    .dma_0_b_valid                                       (dma_bvalid),
    .dma_0_b_bits_id                                     (dma_bid),
    .dma_0_b_bits_resp                                   (dma_bresp),
    .dma_0_ar_ready                                      (dma_arready),
    .dma_0_ar_valid                                      (dma_arvalid),
    .dma_0_ar_bits_id                                    (dma_arid),
    .dma_0_ar_bits_addr                                  (dma_araddr),
    .dma_0_ar_bits_len                                   (dma_arlen),
    .dma_0_ar_bits_size                                  (dma_arsize),
    .dma_0_ar_bits_burst                                 (dma_arburst),
    .dma_0_ar_bits_lock                                  (dma_arlock),
    .dma_0_ar_bits_cache                                 (dma_arcache),
    .dma_0_ar_bits_prot                                  (dma_arprot),
    .dma_0_ar_bits_qos                                   (dma_arqos),
    .dma_0_r_ready                                       (dma_rready),
    .dma_0_r_valid                                       (dma_rvalid),
    .dma_0_r_bits_id                                     (dma_rid),
    .dma_0_r_bits_data                                   (dma_rdata),
    .dma_0_r_bits_resp                                   (dma_rresp),
    .dma_0_r_bits_last                                   (dma_rlast),
    .debug_module_io_resetCtrl_hartResetReq_0
      (_socMisc_debug_module_io_resetCtrl_hartResetReq_0),
    .debug_module_io_resetCtrl_hartIsInReset_0           (_core_with_l2_io_hartIsInReset),
    .debug_module_io_debugIO_clock                       (io_clock),
    .debug_module_io_debugIO_reset                       (_resetGen_o_reset),
    .debug_module_io_debugIO_systemjtag_jtag_TCK         (io_systemjtag_jtag_TCK),
    .debug_module_io_debugIO_systemjtag_jtag_TMS         (io_systemjtag_jtag_TMS),
    .debug_module_io_debugIO_systemjtag_jtag_TDI         (io_systemjtag_jtag_TDI),
    .debug_module_io_debugIO_systemjtag_jtag_TDO_data    (io_systemjtag_jtag_TDO_data),
    .debug_module_io_debugIO_systemjtag_jtag_TDO_driven  (io_systemjtag_jtag_TDO_driven),
    .debug_module_io_debugIO_systemjtag_reset
      (_jtag_reset_sync_resetSync_o_reset),
    .debug_module_io_debugIO_systemjtag_mfr_id           (io_systemjtag_mfr_id),
    .debug_module_io_debugIO_systemjtag_part_number      (io_systemjtag_part_number),
    .debug_module_io_debugIO_systemjtag_version          (io_systemjtag_version),
    .debug_module_io_debugIO_ndreset                     (io_debug_reset),
    .debug_module_io_debugIO_dmactive
      (_socMisc_debug_module_io_debugIO_dmactive),
    .debug_module_io_debugIO_dmactiveAck
      (_socMisc_debug_module_io_debugIO_dmactive),
    .debug_module_io_clock                               (io_clock),
    .debug_module_io_reset                               (_reset_sync_resetSync_o_reset),
    .ext_intrs                                           (io_extIntrs),
    .rtc_clock                                           (io_rtc_clock),
    .pll0_lock                                           (io_pll0_lock),
    .pll0_ctrl_0                                         (io_pll0_ctrl_0),
    .pll0_ctrl_1                                         (io_pll0_ctrl_1),
    .pll0_ctrl_2                                         (io_pll0_ctrl_2),
    .pll0_ctrl_3                                         (io_pll0_ctrl_3),
    .pll0_ctrl_4                                         (io_pll0_ctrl_4),
    .pll0_ctrl_5                                         (io_pll0_ctrl_5),
    .cacheable_check_req_0_bits_addr
      (io_cacheable_check_req_0_bits_addr),
    .cacheable_check_req_1_bits_addr
      (io_cacheable_check_req_1_bits_addr),
    .cacheable_check_resp_0_ld                           (io_cacheable_check_resp_0_ld),
    .cacheable_check_resp_0_st                           (io_cacheable_check_resp_0_st),
    .cacheable_check_resp_0_instr
      (io_cacheable_check_resp_0_instr),
    .cacheable_check_resp_0_mmio                         (io_cacheable_check_resp_0_mmio),
    .cacheable_check_resp_0_atomic
      (io_cacheable_check_resp_0_atomic),
    .cacheable_check_resp_1_ld                           (io_cacheable_check_resp_1_ld),
    .cacheable_check_resp_1_st                           (io_cacheable_check_resp_1_st),
    .cacheable_check_resp_1_instr
      (io_cacheable_check_resp_1_instr),
    .cacheable_check_resp_1_mmio                         (io_cacheable_check_resp_1_mmio),
    .cacheable_check_resp_1_atomic
      (io_cacheable_check_resp_1_atomic),
    .clintTime_valid                                     (_socMisc_clintTime_valid),
    .clintTime_bits                                      (_socMisc_clintTime_bits)
  );
  XSTile core_with_l2 (
    .clock                                                     (io_clock),
    .reset                                                     (_resetGen_1_o_reset),
    .auto_l2top_inner_l2cache_tpmeta_sink_in_valid
      (_broadcast_auto_out_valid),
    .auto_l2top_inner_l2cache_tpmeta_sink_in_bits_hartid
      (_broadcast_auto_out_bits_hartid),
    .auto_l2top_inner_l2cache_tpmeta_sink_in_bits_rawData_0
      (_broadcast_auto_out_bits_rawData_0),
    .auto_l2top_inner_l2cache_tpmeta_sink_in_bits_rawData_1
      (_broadcast_auto_out_bits_rawData_1),
    .auto_l2top_inner_l2cache_tpmeta_sink_in_bits_rawData_2
      (_broadcast_auto_out_bits_rawData_2),
    .auto_l2top_inner_l2cache_tpmeta_source_out_ready
      (_l3cacheOpt_auto_tpmeta_recv_in_ready),
    .auto_l2top_inner_l2cache_tpmeta_source_out_valid
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_valid),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_hartid
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_hartid),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_set
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_set),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_way
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_way),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_wmode
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_wmode),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_0
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_0),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_1
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_1),
    .auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_2
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_2),
    .auto_l2top_inner_beu_int_out_0
      (_core_with_l2_auto_l2top_inner_beu_int_out_0),
    .auto_l2top_inner_nmi_int_in_0                             (nmi_0_0),
    .auto_l2top_inner_nmi_int_in_1                             (nmi_0_1),
    .auto_l2top_inner_plic_int_in_1_0
      (_socMisc_auto_plic_int_out_1_0),
    .auto_l2top_inner_plic_int_in_0_0
      (_socMisc_auto_plic_int_out_0_0),
    .auto_l2top_inner_debug_int_in_0
      (_socMisc_auto_debugModule_debug_dmOuter_dmOuter_int_out_0),
    .auto_l2top_inner_clint_int_in_0
      (_socMisc_auto_clint_int_out_0),
    .auto_l2top_inner_clint_int_in_1
      (_socMisc_auto_clint_int_out_1),
    .auto_l2top_inner_memory_port_out_a_ready
      (_socMisc_auto_buffer_in_a_ready),
    .auto_l2top_inner_memory_port_out_a_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_valid),
    .auto_l2top_inner_memory_port_out_a_bits_opcode
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_opcode),
    .auto_l2top_inner_memory_port_out_a_bits_param
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_param),
    .auto_l2top_inner_memory_port_out_a_bits_size
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_size),
    .auto_l2top_inner_memory_port_out_a_bits_source
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_source),
    .auto_l2top_inner_memory_port_out_a_bits_address
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_address),
    .auto_l2top_inner_memory_port_out_a_bits_user_reqSource
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_user_reqSource),
    .auto_l2top_inner_memory_port_out_a_bits_echo_blockisdirty
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_echo_blockisdirty),
    .auto_l2top_inner_memory_port_out_a_bits_mask
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_mask),
    .auto_l2top_inner_memory_port_out_a_bits_data
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_data),
    .auto_l2top_inner_memory_port_out_a_bits_corrupt
      (_core_with_l2_auto_l2top_inner_memory_port_out_a_bits_corrupt),
    .auto_l2top_inner_memory_port_out_b_ready
      (_core_with_l2_auto_l2top_inner_memory_port_out_b_ready),
    .auto_l2top_inner_memory_port_out_b_valid
      (_socMisc_auto_buffer_in_b_valid),
    .auto_l2top_inner_memory_port_out_b_bits_opcode
      (_socMisc_auto_buffer_in_b_bits_opcode),
    .auto_l2top_inner_memory_port_out_b_bits_param
      (_socMisc_auto_buffer_in_b_bits_param),
    .auto_l2top_inner_memory_port_out_b_bits_size
      (_socMisc_auto_buffer_in_b_bits_size),
    .auto_l2top_inner_memory_port_out_b_bits_address
      (_socMisc_auto_buffer_in_b_bits_address),
    .auto_l2top_inner_memory_port_out_b_bits_mask
      (_socMisc_auto_buffer_in_b_bits_mask),
    .auto_l2top_inner_memory_port_out_b_bits_data
      (_socMisc_auto_buffer_in_b_bits_data),
    .auto_l2top_inner_memory_port_out_b_bits_corrupt
      (_socMisc_auto_buffer_in_b_bits_corrupt),
    .auto_l2top_inner_memory_port_out_c_ready
      (_socMisc_auto_buffer_in_c_ready),
    .auto_l2top_inner_memory_port_out_c_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_valid),
    .auto_l2top_inner_memory_port_out_c_bits_opcode
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_opcode),
    .auto_l2top_inner_memory_port_out_c_bits_param
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_param),
    .auto_l2top_inner_memory_port_out_c_bits_size
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_size),
    .auto_l2top_inner_memory_port_out_c_bits_source
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_source),
    .auto_l2top_inner_memory_port_out_c_bits_address
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_address),
    .auto_l2top_inner_memory_port_out_c_bits_user_reqSource
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_user_reqSource),
    .auto_l2top_inner_memory_port_out_c_bits_echo_blockisdirty
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_echo_blockisdirty),
    .auto_l2top_inner_memory_port_out_c_bits_data
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_data),
    .auto_l2top_inner_memory_port_out_c_bits_corrupt
      (_core_with_l2_auto_l2top_inner_memory_port_out_c_bits_corrupt),
    .auto_l2top_inner_memory_port_out_d_ready
      (_core_with_l2_auto_l2top_inner_memory_port_out_d_ready),
    .auto_l2top_inner_memory_port_out_d_valid
      (_socMisc_auto_buffer_in_d_valid),
    .auto_l2top_inner_memory_port_out_d_bits_opcode
      (_socMisc_auto_buffer_in_d_bits_opcode),
    .auto_l2top_inner_memory_port_out_d_bits_param
      (_socMisc_auto_buffer_in_d_bits_param),
    .auto_l2top_inner_memory_port_out_d_bits_size
      (_socMisc_auto_buffer_in_d_bits_size),
    .auto_l2top_inner_memory_port_out_d_bits_source
      (_socMisc_auto_buffer_in_d_bits_source),
    .auto_l2top_inner_memory_port_out_d_bits_sink
      (_socMisc_auto_buffer_in_d_bits_sink),
    .auto_l2top_inner_memory_port_out_d_bits_denied
      (_socMisc_auto_buffer_in_d_bits_denied),
    .auto_l2top_inner_memory_port_out_d_bits_echo_blockisdirty
      (_socMisc_auto_buffer_in_d_bits_echo_blockisdirty),
    .auto_l2top_inner_memory_port_out_d_bits_data
      (_socMisc_auto_buffer_in_d_bits_data),
    .auto_l2top_inner_memory_port_out_d_bits_corrupt
      (_socMisc_auto_buffer_in_d_bits_corrupt),
    .auto_l2top_inner_memory_port_out_e_ready
      (_socMisc_auto_buffer_in_e_ready),
    .auto_l2top_inner_memory_port_out_e_valid
      (_core_with_l2_auto_l2top_inner_memory_port_out_e_valid),
    .auto_l2top_inner_memory_port_out_e_bits_sink
      (_core_with_l2_auto_l2top_inner_memory_port_out_e_bits_sink),
    .auto_l2top_inner_mmio_port_out_a_ready
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_a_ready),
    .auto_l2top_inner_mmio_port_out_a_valid
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_valid),
    .auto_l2top_inner_mmio_port_out_a_bits_opcode
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_opcode),
    .auto_l2top_inner_mmio_port_out_a_bits_param
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_param),
    .auto_l2top_inner_mmio_port_out_a_bits_size
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_size),
    .auto_l2top_inner_mmio_port_out_a_bits_source
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_source),
    .auto_l2top_inner_mmio_port_out_a_bits_address
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_address),
    .auto_l2top_inner_mmio_port_out_a_bits_mask
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_mask),
    .auto_l2top_inner_mmio_port_out_a_bits_data
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_data),
    .auto_l2top_inner_mmio_port_out_a_bits_corrupt
      (_core_with_l2_auto_l2top_inner_mmio_port_out_a_bits_corrupt),
    .auto_l2top_inner_mmio_port_out_d_ready
      (_core_with_l2_auto_l2top_inner_mmio_port_out_d_ready),
    .auto_l2top_inner_mmio_port_out_d_valid
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_valid),
    .auto_l2top_inner_mmio_port_out_d_bits_opcode
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_opcode),
    .auto_l2top_inner_mmio_port_out_d_bits_param
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_param),
    .auto_l2top_inner_mmio_port_out_d_bits_size
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_size),
    .auto_l2top_inner_mmio_port_out_d_bits_source
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_source),
    .auto_l2top_inner_mmio_port_out_d_bits_sink
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_sink),
    .auto_l2top_inner_mmio_port_out_d_bits_denied
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_denied),
    .auto_l2top_inner_mmio_port_out_d_bits_data
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_data),
    .auto_l2top_inner_mmio_port_out_d_bits_corrupt
      (_socMisc_auto_L2_to_L3_peripheral_buffer_1_in_d_bits_corrupt),
    .auto_core_memBlock_inner_l3_pf_sender_out_addr
      (_core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr),
    .auto_core_memBlock_inner_l3_pf_sender_out_addr_valid
      (_core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr_valid),
    .io_hartId                                                 (6'h0),
    .io_msiInfo_valid                                          (1'h0),
    .io_msiInfo_bits_info                                      (17'h0),
    .io_reset_vector                                           (io_riscv_rst_vec_0),
    .io_cpu_halt                                               (io_riscv_halt_0),
    .io_cpu_poff                                               (/* unused */),
    .io_cpu_crtical_error
      (io_riscv_critical_error_0),
    .io_hartIsInReset
      (_core_with_l2_io_hartIsInReset),
    .io_traceCoreInterface_fromEncoder_enable
      (io_traceCoreInterface_0_fromEncoder_enable),
    .io_traceCoreInterface_fromEncoder_stall
      (io_traceCoreInterface_0_fromEncoder_stall),
    .io_traceCoreInterface_toEncoder_priv
      (io_traceCoreInterface_0_toEncoder_priv),
    .io_traceCoreInterface_toEncoder_trap_cause
      (io_traceCoreInterface_0_toEncoder_cause),
    .io_traceCoreInterface_toEncoder_trap_tval
      (io_traceCoreInterface_0_toEncoder_tval),
    .io_traceCoreInterface_toEncoder_groups_0_bits_iaddr
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iaddr),
    .io_traceCoreInterface_toEncoder_groups_0_bits_itype
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_itype),
    .io_traceCoreInterface_toEncoder_groups_0_bits_iretire
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iretire),
    .io_traceCoreInterface_toEncoder_groups_0_bits_ilastsize
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_ilastsize),
    .io_traceCoreInterface_toEncoder_groups_1_bits_iaddr
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iaddr),
    .io_traceCoreInterface_toEncoder_groups_1_bits_itype
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_itype),
    .io_traceCoreInterface_toEncoder_groups_1_bits_iretire
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iretire),
    .io_traceCoreInterface_toEncoder_groups_1_bits_ilastsize
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_ilastsize),
    .io_traceCoreInterface_toEncoder_groups_2_bits_iaddr
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iaddr),
    .io_traceCoreInterface_toEncoder_groups_2_bits_itype
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_itype),
    .io_traceCoreInterface_toEncoder_groups_2_bits_iretire
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iretire),
    .io_traceCoreInterface_toEncoder_groups_2_bits_ilastsize
      (_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_ilastsize),
    .io_l3Miss                                                 (_l3cacheOpt_io_l3Miss),
    .io_clintTime_valid                                        (_socMisc_clintTime_valid),
    .io_clintTime_bits                                         (_socMisc_clintTime_bits)
  );
  HuanCun l3cacheOpt (
    .clock                                (io_clock),
    .reset                                (_resetGen_o_reset),
    .auto_ctrl_unit_int_out_0             (_l3cacheOpt_auto_ctrl_unit_int_out_0),
    .auto_ctrl_unit_ctl_in_a_ready        (_l3cacheOpt_auto_ctrl_unit_ctl_in_a_ready),
    .auto_ctrl_unit_ctl_in_a_valid        (_socMisc_auto_xbar_out_0_a_valid),
    .auto_ctrl_unit_ctl_in_a_bits_opcode  (_socMisc_auto_xbar_out_0_a_bits_opcode),
    .auto_ctrl_unit_ctl_in_a_bits_size    (_socMisc_auto_xbar_out_0_a_bits_size),
    .auto_ctrl_unit_ctl_in_a_bits_source  (_socMisc_auto_xbar_out_0_a_bits_source),
    .auto_ctrl_unit_ctl_in_a_bits_address (_socMisc_auto_xbar_out_0_a_bits_address),
    .auto_ctrl_unit_ctl_in_a_bits_mask    (_socMisc_auto_xbar_out_0_a_bits_mask),
    .auto_ctrl_unit_ctl_in_a_bits_data    (_socMisc_auto_xbar_out_0_a_bits_data),
    .auto_ctrl_unit_ctl_in_d_ready        (_socMisc_auto_xbar_out_0_d_ready),
    .auto_ctrl_unit_ctl_in_d_valid        (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_valid),
    .auto_ctrl_unit_ctl_in_d_bits_opcode
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_opcode),
    .auto_ctrl_unit_ctl_in_d_bits_size    (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_size),
    .auto_ctrl_unit_ctl_in_d_bits_source
      (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_source),
    .auto_ctrl_unit_ctl_in_d_bits_data    (_l3cacheOpt_auto_ctrl_unit_ctl_in_d_bits_data),
    .auto_tpmeta_send_out_valid           (_l3cacheOpt_auto_tpmeta_send_out_valid),
    .auto_tpmeta_send_out_bits_hartid     (_l3cacheOpt_auto_tpmeta_send_out_bits_hartid),
    .auto_tpmeta_send_out_bits_rawData_0
      (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_0),
    .auto_tpmeta_send_out_bits_rawData_1
      (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_1),
    .auto_tpmeta_send_out_bits_rawData_2
      (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_2),
    .auto_tpmeta_recv_in_ready            (_l3cacheOpt_auto_tpmeta_recv_in_ready),
    .auto_tpmeta_recv_in_valid
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_valid),
    .auto_tpmeta_recv_in_bits_hartid
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_hartid),
    .auto_tpmeta_recv_in_bits_set
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_set),
    .auto_tpmeta_recv_in_bits_way
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_way),
    .auto_tpmeta_recv_in_bits_wmode
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_wmode),
    .auto_tpmeta_recv_in_bits_rawData_0
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_0),
    .auto_tpmeta_recv_in_bits_rawData_1
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_1),
    .auto_tpmeta_recv_in_bits_rawData_2
      (_core_with_l2_auto_l2top_inner_l2cache_tpmeta_source_out_bits_rawData_2),
    .auto_pf_recv_in_addr
      (_core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr),
    .auto_pf_recv_in_addr_valid
      (_core_with_l2_auto_core_memBlock_inner_l3_pf_sender_out_addr_valid),
    .auto_in_a_ready                      (_l3cacheOpt_auto_in_a_ready),
    .auto_in_a_valid                      (_socMisc_auto_xbar_out_1_a_valid),
    .auto_in_a_bits_opcode                (_socMisc_auto_xbar_out_1_a_bits_opcode),
    .auto_in_a_bits_param                 (_socMisc_auto_xbar_out_1_a_bits_param),
    .auto_in_a_bits_size                  (_socMisc_auto_xbar_out_1_a_bits_size),
    .auto_in_a_bits_source                (_socMisc_auto_xbar_out_1_a_bits_source),
    .auto_in_a_bits_address               (_socMisc_auto_xbar_out_1_a_bits_address),
    .auto_in_a_bits_user_reqSource
      (_socMisc_auto_xbar_out_1_a_bits_user_reqSource),
    .auto_in_a_bits_mask                  (_socMisc_auto_xbar_out_1_a_bits_mask),
    .auto_in_a_bits_data                  (_socMisc_auto_xbar_out_1_a_bits_data),
    .auto_in_a_bits_corrupt               (_socMisc_auto_xbar_out_1_a_bits_corrupt),
    .auto_in_b_ready                      (_socMisc_auto_xbar_out_1_b_ready),
    .auto_in_b_valid                      (_l3cacheOpt_auto_in_b_valid),
    .auto_in_b_bits_param                 (_l3cacheOpt_auto_in_b_bits_param),
    .auto_in_b_bits_address               (_l3cacheOpt_auto_in_b_bits_address),
    .auto_in_b_bits_data                  (_l3cacheOpt_auto_in_b_bits_data),
    .auto_in_c_ready                      (_l3cacheOpt_auto_in_c_ready),
    .auto_in_c_valid                      (_socMisc_auto_xbar_out_1_c_valid),
    .auto_in_c_bits_opcode                (_socMisc_auto_xbar_out_1_c_bits_opcode),
    .auto_in_c_bits_param                 (_socMisc_auto_xbar_out_1_c_bits_param),
    .auto_in_c_bits_size                  (_socMisc_auto_xbar_out_1_c_bits_size),
    .auto_in_c_bits_source                (_socMisc_auto_xbar_out_1_c_bits_source),
    .auto_in_c_bits_address               (_socMisc_auto_xbar_out_1_c_bits_address),
    .auto_in_c_bits_echo_blockisdirty
      (_socMisc_auto_xbar_out_1_c_bits_echo_blockisdirty),
    .auto_in_c_bits_data                  (_socMisc_auto_xbar_out_1_c_bits_data),
    .auto_in_d_ready                      (_socMisc_auto_xbar_out_1_d_ready),
    .auto_in_d_valid                      (_l3cacheOpt_auto_in_d_valid),
    .auto_in_d_bits_opcode                (_l3cacheOpt_auto_in_d_bits_opcode),
    .auto_in_d_bits_param                 (_l3cacheOpt_auto_in_d_bits_param),
    .auto_in_d_bits_size                  (_l3cacheOpt_auto_in_d_bits_size),
    .auto_in_d_bits_source                (_l3cacheOpt_auto_in_d_bits_source),
    .auto_in_d_bits_sink                  (_l3cacheOpt_auto_in_d_bits_sink),
    .auto_in_d_bits_denied                (_l3cacheOpt_auto_in_d_bits_denied),
    .auto_in_d_bits_echo_blockisdirty     (_l3cacheOpt_auto_in_d_bits_echo_blockisdirty),
    .auto_in_d_bits_data                  (_l3cacheOpt_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt               (_l3cacheOpt_auto_in_d_bits_corrupt),
    .auto_in_e_valid                      (_socMisc_auto_xbar_out_1_e_valid),
    .auto_in_e_bits_sink                  (_socMisc_auto_xbar_out_1_e_bits_sink),
    .auto_out_a_ready                     (_socMisc_auto_binder_in_a_ready),
    .auto_out_a_valid                     (_l3cacheOpt_auto_out_a_valid),
    .auto_out_a_bits_opcode               (_l3cacheOpt_auto_out_a_bits_opcode),
    .auto_out_a_bits_param                (_l3cacheOpt_auto_out_a_bits_param),
    .auto_out_a_bits_size                 (_l3cacheOpt_auto_out_a_bits_size),
    .auto_out_a_bits_source               (_l3cacheOpt_auto_out_a_bits_source),
    .auto_out_a_bits_address              (_l3cacheOpt_auto_out_a_bits_address),
    .auto_out_a_bits_mask                 (_l3cacheOpt_auto_out_a_bits_mask),
    .auto_out_a_bits_data                 (_l3cacheOpt_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt              (_l3cacheOpt_auto_out_a_bits_corrupt),
    .auto_out_c_ready                     (_socMisc_auto_binder_in_c_ready),
    .auto_out_c_valid                     (_l3cacheOpt_auto_out_c_valid),
    .auto_out_c_bits_opcode               (_l3cacheOpt_auto_out_c_bits_opcode),
    .auto_out_c_bits_size                 (_l3cacheOpt_auto_out_c_bits_size),
    .auto_out_c_bits_source               (_l3cacheOpt_auto_out_c_bits_source),
    .auto_out_c_bits_address              (_l3cacheOpt_auto_out_c_bits_address),
    .auto_out_c_bits_data                 (_l3cacheOpt_auto_out_c_bits_data),
    .auto_out_c_bits_corrupt              (_l3cacheOpt_auto_out_c_bits_corrupt),
    .auto_out_d_ready                     (_l3cacheOpt_auto_out_d_ready),
    .auto_out_d_valid                     (_socMisc_auto_binder_in_d_valid),
    .auto_out_d_bits_opcode               (_socMisc_auto_binder_in_d_bits_opcode),
    .auto_out_d_bits_param                (_socMisc_auto_binder_in_d_bits_param),
    .auto_out_d_bits_size                 (_socMisc_auto_binder_in_d_bits_size),
    .auto_out_d_bits_source               (_socMisc_auto_binder_in_d_bits_source),
    .auto_out_d_bits_sink                 (_socMisc_auto_binder_in_d_bits_sink),
    .auto_out_d_bits_denied               (_socMisc_auto_binder_in_d_bits_denied),
    .auto_out_d_bits_data                 (_socMisc_auto_binder_in_d_bits_data),
    .auto_out_d_bits_corrupt              (_socMisc_auto_binder_in_d_bits_corrupt),
    .auto_out_e_valid                     (_l3cacheOpt_auto_out_e_valid),
    .auto_out_e_bits_sink                 (_l3cacheOpt_auto_out_e_bits_sink),
    .io_l3Miss                            (_l3cacheOpt_io_l3Miss)
  );
  IntBuffer intBuffer (
    .clock      (io_clock),
    .reset      (_reset_sync_resetSync_o_reset),
    .auto_in_0  (_core_with_l2_auto_l2top_inner_beu_int_out_0),
    .auto_out_0 (_intBuffer_auto_out_0)
  );
  IntBuffer intBuffer_1 (
    .clock      (io_clock),
    .reset      (_reset_sync_resetSync_o_reset),
    .auto_in_0  (_l3cacheOpt_auto_ctrl_unit_int_out_0),
    .auto_out_0 (_intBuffer_1_auto_out_0)
  );
  ValidIOBroadcast broadcast (
    .auto_in_valid           (_l3cacheOpt_auto_tpmeta_send_out_valid),
    .auto_in_bits_hartid     (_l3cacheOpt_auto_tpmeta_send_out_bits_hartid),
    .auto_in_bits_rawData_0  (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_0),
    .auto_in_bits_rawData_1  (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_1),
    .auto_in_bits_rawData_2  (_l3cacheOpt_auto_tpmeta_send_out_bits_rawData_2),
    .auto_out_valid          (_broadcast_auto_out_valid),
    .auto_out_bits_hartid    (_broadcast_auto_out_bits_hartid),
    .auto_out_bits_rawData_0 (_broadcast_auto_out_bits_rawData_0),
    .auto_out_bits_rawData_1 (_broadcast_auto_out_bits_rawData_1),
    .auto_out_bits_rawData_2 (_broadcast_auto_out_bits_rawData_2)
  );
  ResetGen reset_sync_resetSync (
    .clock   (io_clock),
    .reset   (io_reset),
    .o_reset (_reset_sync_resetSync_o_reset)
  );
  ResetGen jtag_reset_sync_resetSync (
    .clock   (io_systemjtag_jtag_TCK),
    .reset   (io_systemjtag_reset),
    .o_reset (_jtag_reset_sync_resetSync_o_reset)
  );
  ResetGen resetGen (
    .clock   (io_clock),
    .reset   (_reset_sync_resetSync_o_reset),
    .o_reset (_resetGen_o_reset)
  );
  ResetGen resetGen_1 (
    .clock   (io_clock),
    .reset   (_resetGen_o_reset | _socMisc_debug_module_io_resetCtrl_hartResetReq_0),
    .o_reset (_resetGen_1_o_reset)
  );
  assign io_traceCoreInterface_0_toEncoder_iaddr =
    {_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iaddr,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iaddr,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iaddr};
  assign io_traceCoreInterface_0_toEncoder_itype =
    {_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_itype,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_itype,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_itype};
  assign io_traceCoreInterface_0_toEncoder_iretire =
    {_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_iretire,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_iretire,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_iretire};
  assign io_traceCoreInterface_0_toEncoder_ilastsize =
    {_core_with_l2_io_traceCoreInterface_toEncoder_groups_2_bits_ilastsize,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_1_bits_ilastsize,
     _core_with_l2_io_traceCoreInterface_toEncoder_groups_0_bits_ilastsize};
endmodule

